module tb_execute();
    logic		clk;
    logic 		fowarded_data;
    logic [24:0]	instructionID;
    logic [127:0]	rs1, rs2, rs3; 
    logic [127:0]	ALUOut;
    logic [24:0]	instructionWB;
    logic [31:0]	word1, word2, word3, word4;
    logic [15:0]	hw1, hw2, hw3, hw4, hw5, hw6, hw7, hw8;
    logic [63:0]	long1, long2;

    execute U0(
	.rs1 (rs1),
	.rs2 (rs2),
	.rs3 (rs3),
	.fowarded_data (fowarded_data),
	.instructionID (instructionID),
	.ALUOut (ALUOut),
	.instructionWB (instructionWB));


    initial begin
	clk = 0;
	/*//A
	instructionID = 25'b1100000001000000000000000;	//5 + 6 4x
	rs1 = 5;
	rs2 = 6;
	rs1[63:32] = -5;
	rs1[95:64] = 20000;
	rs1[127:96] = -20000;
	rs2[63:32] = -6;
	rs2[95:64] = 20000;
	rs2[127:96] = -20000;*/
	
	//AH
/*	instructionID = 25'b1100000010000000000000000;	//5 + 6 4x
	rs1[15:0] = -5;
	rs1[31:16] = 20000;
	rs1[47:32] = -20000;
	rs1[63:48] = -6;
	rs1[79:64] = 20000;
	rs1[95:80] = -20000;
	rs1[111:96] = -5;
	rs1[127:112] = 20000;

	rs2[15:0] = -5;
	rs2[31:16] = 20000;
	rs2[47:32] = -20000;
	rs2[63:48] = -6;
	rs2[79:64] = 20000;
	rs2[95:80] = -20000;
	rs2[111:96] = -5;
	rs2[127:112] = 20000;*/


	//MPYU cant overflow
/*	instructionID = 25'b1100001010000000000000000;	
	rs1[15:0] = 1;
	rs1[31:16] = 0;
	rs1[47:32] = 200;
	rs1[63:48] = 0;
	rs1[79:64] = 40000;
	rs1[95:80] = 0;
	rs1[111:96] = 3;
	rs1[127:112] = 1;

	rs2[15:0] = 1;
	rs2[31:16] = 0;
	rs2[47:32] = 200;
	rs2[63:48] = 0;
	rs2[79:64] = 40000;//overflow
	rs2[95:80] = 0;
	rs2[111:96] = 0;
	rs2[127:112] = 1;*/

	//OR
/*	instructionID = 25'b1100001011000000000000000;	
	rs1[63:0] = 64'hFFFFFFFF00000000;
	rs1[127:64] = 64'hFFFFFFFFFFFFFFFF;

	rs2[63:0] = 64'hFFFFFFFF00000000;
	rs2[127:64] = 64'h0000000000000000;*/

	//POPCNT
/*	instructionID = 25'b1100001100000000000000000;	
	rs1[15:0] = 1;
	rs1[31:16] = 3;
	rs1[47:32] = 7;
	rs1[63:48] = 15;
	rs1[79:64] = 31;
	rs1[95:80] = 63;
	rs1[111:96] = 127;
	rs1[127:112] = 255;

	rs2[15:0] = 0;
	rs2[31:16] = 0;
	rs2[47:32] = 0;
	rs2[63:48] = 0;
	rs2[79:64] = 0;//overflow
	rs2[95:80] = 0;
	rs2[111:96] = 0;
	rs2[127:112] = 0;*/

	//ROT
/*	instructionID = 25'b1100001101000000000000000;	
	rs1[127:0] = 15;

	rs2[127:0] = 1;
*/

	//ROTW
/*	instructionID = 25'b1100001110000000000000000;	
	//rs1[15:0] = 15;
	rs1[31:0] = 15;
	//rs1[47:32] = 15;
	rs1[63:32] = 15;
	//rs1[79:64] = 15;
	rs1[95:64] = 15;
	//rs1[111:96] = 15;
	rs1[127:96] = 15;

	//rs1[15:0] = 15;
	rs2[31:0] = 1;
	//rs1[47:32] = 15;
	rs2[63:32] = 2;
	//rs1[79:64] = 15;
	rs2[95:64] = 3;
	//rs1[111:96] = 15;
	rs2[127:96] = 4;*/

	//SHLHI
/*	instructionID = 25'b1100001111000000000000000;	
	rs1[15:0] = 15;
	rs1[31:16] = 15;
	rs1[47:32] = 15;
	rs1[63:48] = 15;
	rs1[79:64] = 15;
	rs1[95:80] = 15;
	rs1[111:96] = 15;
	rs1[127:112] = 15;

	rs2[15:0] = 1;
	rs2[31:16] = 2;
	rs2[47:32] = 3;
	rs2[63:48] = 4;
	rs2[79:64] = 5;
	rs2[95:80] = 6;
	rs2[111:96] = 7;
	rs2[127:112] = 8;*/

	//SFH
/*	instructionID = 25'b1100010000000000000000000;	
	rs1[15:0] = 15;
	rs1[31:16] = 15;
	rs1[47:32] = 15;
	rs1[63:48] = 15;
	rs1[79:64] = 15;
	rs1[95:80] = 15;
	rs1[111:96] = 7;
	rs1[127:112] = 7;

	rs2[15:0] = 1;
	rs2[31:16] = 2;
	rs2[47:32] = 3;
	rs2[63:48] = 4;
	rs2[79:64] = 5;
	rs2[95:80] = 6;
	rs2[111:96] = 7;
	rs2[127:112] = 8;*/

	//SFW
/*	instructionID = 25'b1100010001000000000000000;	
	//rs1[15:0] = 15;
	rs1[31:0] = 15;
	//rs1[47:32] = 15;
	rs1[63:32] = 15;
	//rs1[79:64] = 15;
	rs1[95:64] = 15;
	//rs1[111:96] = 7;
	rs1[127:96] = 7;

	//rs2[15:0] = 1;
	rs2[31:0] = 1;
	//rs2[47:32] = 3;
	rs2[63:32] = 2;
	//rs2[79:64] = 5;
	rs2[95:64] = 15;
	//rs2[111:96] = 7;
	rs2[127:96] = 8;*/

	//SFHS
/*	instructionID = 25'b1100010010000000000000000;	
	rs1[15:0] = 15;
	rs1[31:16] = 15;
	rs1[47:32] = -1;
	rs1[63:48] = -2;
	rs1[79:64] = 15;
	rs1[95:80] = 15;
	rs1[111:96] = 7;
	rs1[127:112] = -32767;

	rs2[15:0] = 16;
	rs2[31:16] = 14;
	rs2[47:32] = -2;
	rs2[63:48] = -1;
	rs2[79:64] = 5;
	rs2[95:80] = 6;
	rs2[111:96] = 7;
	rs2[127:112] = 8;*/

	//XOR
/*	instructionID = 25'b1100010011000000000000000;	
	rs1[63:0] = 64'hFFFFFFFF00000000;
	rs1[127:64] = 64'hFFFFFFFFFFFFFFFF;

	rs2[63:0] = 64'hFFFFFFFF00000000;
	rs2[127:64] = 64'h0000000000000000;*/

	//A
/*	instructionID = 25'b1100000001000000000000000;	
	//rs1[15:0] = 15;
	rs1[31:0] = 1;
	//rs1[47:32] = 15;
	rs1[63:32] = 2;
	//rs1[79:64] = 15;
	rs1[95:64] = 3;
	//rs1[111:96] = 7;
	rs1[127:96] = 33'd4294967296;

	//rs2[15:0] = 1;
	rs2[31:0] = 1;
	//rs2[47:32] = 3;
	rs2[63:32] = 2;
	//rs2[79:64] = 5;
	rs2[95:64] = 3;
	//rs2[111:96] = 7;
	rs2[127:96] = 2;*/

	//AH
/*	instructionID = 25'b1100000010000000000000000;	
	rs1[15:0] = 15;
	rs1[31:16] = 15;
	rs1[47:32] = 15;
	rs1[63:48] = 15;
	rs1[79:64] = 15;
	rs1[95:80] = 15;
	rs1[111:96] = 15;
	rs1[127:112] = 17'd65535;

	rs2[15:0] = 1;
	rs2[31:16] = 2;
	rs2[47:32] = 3;
	rs2[63:48] = 4;
	rs2[79:64] = 5;
	rs2[95:80] = 6;
	rs2[111:96] = 7;
	rs2[127:112] = 8;*/

	//AHS
/*	instructionID = 25'b1100000011000000000000000;	
	rs1[15:0] = 15;
	rs1[31:16] = 15;
	rs1[47:32] = 15;
	rs1[63:48] = 15;
	rs1[79:64] = 15;
	rs1[95:80] = 15;
	rs1[111:96] = 15;
	rs1[127:112] = 17'd32767;

	rs2[15:0] = 1;
	rs2[31:16] = 2;
	rs2[47:32] = 3;
	rs2[63:48] = 4;
	rs2[79:64] = 5;
	rs2[95:80] = 6;
	rs2[111:96] = 7;
	rs2[127:112] = 8;*/

	//AND
/*	instructionID = 25'b1100000100000000000000000;	
	rs1[63:0] = 64'hFFFFFFFF00000000;
	rs1[127:64] = 64'hFFFFFFFFFFFFFFFF;

	rs2[63:0] = 64'hFFFFFFFF00000000;
	rs2[127:64] = 64'h0000000000000000;*/

	//BCW
/*	instructionID = 25'b1100000101000000000000000;	
	rs1[63:0] = 64'h00000000FFFFFFFE;
	rs1[127:64] = 64'h0000000000000000;

	rs2[63:0] = 64'h0000000000000000;
	rs2[127:64] = 64'h0000000000000000;*/

	//CLZ
/*	instructionID = 25'b1100000110000000000000000;	
	rs1[63:0] = 64'h000000000FFFFFFE;
	rs1[127:64] = 64'h0000000000000001;

	rs2[63:0] = 64'h0000000000000000;
	rs2[127:64] = 64'h0000000000000000;*/


	//MAX
	/*instructionID = 25'b1100000111000000000000000;	
	//rs1[15:0] = 15;
	rs1[31:0] = -1;
	//rs1[47:32] = 15;
	rs1[63:32] = -2;
	//rs1[79:64] = 15;
	rs1[95:64] = -100;
	//rs1[111:96] = 7;
	rs1[127:96] = 0;

	//rs2[15:0] = 1;
	rs2[31:0] = -8;
	//rs2[47:32] = 3;
	rs2[63:32] = -8;
	//rs2[79:64] = 5;
	rs2[95:64] = -3;
	//rs2[111:96] = 7;
	rs2[127:96] = -33'd4294967296;*/

	//MIN
/*	instructionID = 25'b1100001000000000000000000;	
	//rs1[15:0] = 15;
	rs1[31:0] = 1;
	//rs1[47:32] = 15;
	rs1[63:32] = 2;
	//rs1[79:64] = 15;
	rs1[95:64] = 100;
	//rs1[111:96] = 7;
	rs1[127:96] = 0;

	//rs2[15:0] = 1;
	rs2[31:0] = 8;
	//rs2[47:32] = 3;
	rs2[63:32] = 8;
	//rs2[79:64] = 5;
	rs2[95:64] = 3;
	//rs2[111:96] = 7;
	rs2[127:96] = -32'd2147483648;*/

	//MSGN
	instructionID = 25'b1100001001000000000000000;	
	//rs1[15:0] = 15;
	rs1[31:0] = -32'd2147483648;
	//rs1[47:32] = 15;
	rs1[63:32] = 0;
	//rs1[79:64] = 15;
	rs1[95:64] = 100;
	//rs1[111:96] = 7;
	rs1[127:96] = 100;

	rs2[31:0]=0;
	rs2[63]=1;
	rs2[95]=1;
	rs2[127]=0;


    end

    always begin
	#1 clk = !clk;
	word1 = ALUOut[31:0];
	word2 = ALUOut[63:32];
	word3 = ALUOut[95:64];
	word4 = ALUOut[127:96];
	hw1 = ALUOut[15:0];
	hw2 = ALUOut[31:16];
	hw3 = ALUOut[47:32];
	hw4 = ALUOut[63:48];
	hw5 = ALUOut[79:64];
	hw6 = ALUOut[95:80];
	hw7 = ALUOut[111:96];
	hw8 = ALUOut[127:112];
	long1 = ALUOut[63:0];
	long2 = ALUOut[127:64];
    end

    initial begin
	#100;
	$finish;
    end

endmodule
		







